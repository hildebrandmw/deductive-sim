module test_not(N1, N2);

input N1;
output N2;

not INV1_1 (N2, N1);

endmodule
