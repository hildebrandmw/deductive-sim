module test_or(N3, N2, N1);

input N1,N2;
output N3;


or OR2_1 (N3, N2, N1);
endmodule
