module test_nand(N3, N2, N1);

input N1,N2;
output N3;


nand NAND2_1 (N3, N2, N1);
endmodule
