module c7552_tb();
parameter INPUT_WIDTH = 207;
parameter OUTPUT_WIDTH = 108;
parameter NUMBER_OF_TESTS = 10000;
string INPUT_FILE = "input_vectors/c7552.txt";
string OUTPUT_FILE = "output_vectors/c7552.txt";

reg   [INPUT_WIDTH-1:0] in;
wire  [OUTPUT_WIDTH-1:0] out;

reg [INPUT_WIDTH-1:0] memory [NUMBER_OF_TESTS-1:0];
integer i,f;

c7552 UUT (.N1(in[0]), .N5(in[1]), .N9(in[2]), .N12(in[3]), 
.N15(in[4]), .N18(in[5]), .N23(in[6]), .N26(in[7]), 
.N29(in[8]), .N32(in[9]), .N35(in[10]), .N38(in[11]), 
.N41(in[12]), .N44(in[13]), .N47(in[14]), .N50(in[15]), 
.N53(in[16]), .N54(in[17]), .N55(in[18]), .N56(in[19]), 
.N57(in[20]), .N58(in[21]), .N59(in[22]), .N60(in[23]), 
.N61(in[24]), .N62(in[25]), .N63(in[26]), .N64(in[27]), 
.N65(in[28]), .N66(in[29]), .N69(in[30]), .N70(in[31]), 
.N73(in[32]), .N74(in[33]), .N75(in[34]), .N76(in[35]), 
.N77(in[36]), .N78(in[37]), .N79(in[38]), .N80(in[39]), 
.N81(in[40]), .N82(in[41]), .N83(in[42]), .N84(in[43]), 
.N85(in[44]), .N86(in[45]), .N87(in[46]), .N88(in[47]), 
.N89(in[48]), .N94(in[49]), .N97(in[50]), .N100(in[51]), 
.N103(in[52]), .N106(in[53]), .N109(in[54]), .N110(in[55]), 
.N111(in[56]), .N112(in[57]), .N113(in[58]), .N114(in[59]), 
.N115(in[60]), .N118(in[61]), .N121(in[62]), .N124(in[63]), 
.N127(in[64]), .N130(in[65]), .N133(in[66]), .N134(in[67]), 
.N135(in[68]), .N138(in[69]), .N141(in[70]), .N144(in[71]), 
.N147(in[72]), .N150(in[73]), .N151(in[74]), .N152(in[75]), 
.N153(in[76]), .N154(in[77]), .N155(in[78]), .N156(in[79]), 
.N157(in[80]), .N158(in[81]), .N159(in[82]), .N160(in[83]), 
.N161(in[84]), .N162(in[85]), .N163(in[86]), .N164(in[87]), 
.N165(in[88]), .N166(in[89]), .N167(in[90]), .N168(in[91]), 
.N169(in[92]), .N170(in[93]), .N171(in[94]), .N172(in[95]), 
.N173(in[96]), .N174(in[97]), .N175(in[98]), .N176(in[99]), 
.N177(in[100]), .N178(in[101]), .N179(in[102]), .N180(in[103]), 
.N181(in[104]), .N182(in[105]), .N183(in[106]), .N184(in[107]), 
.N185(in[108]), .N186(in[109]), .N187(in[110]), .N188(in[111]), 
.N189(in[112]), .N190(in[113]), .N191(in[114]), .N192(in[115]), 
.N193(in[116]), .N194(in[117]), .N195(in[118]), .N196(in[119]), 
.N197(in[120]), .N198(in[121]), .N199(in[122]), .N200(in[123]), 
.N201(in[124]), .N202(in[125]), .N203(in[126]), .N204(in[127]), 
.N205(in[128]), .N206(in[129]), .N207(in[130]), .N208(in[131]), 
.N209(in[132]), .N210(in[133]), .N211(in[134]), .N212(in[135]), 
.N213(in[136]), .N214(in[137]), .N215(in[138]), .N216(in[139]), 
.N217(in[140]), .N218(in[141]), .N219(in[142]), .N220(in[143]), 
.N221(in[144]), .N222(in[145]), .N223(in[146]), .N224(in[147]), 
.N225(in[148]), .N226(in[149]), .N227(in[150]), .N228(in[151]), 
.N229(in[152]), .N230(in[153]), .N231(in[154]), .N232(in[155]), 
.N233(in[156]), .N234(in[157]), .N235(in[158]), .N236(in[159]), 
.N237(in[160]), .N238(in[161]), .N239(in[162]), .N240(in[163]), 
.N242(in[164]), .N245(in[165]), .N248(in[166]), .N251(in[167]), 
.N254(in[168]), .N257(in[169]), .N260(in[170]), .N263(in[171]), 
.N267(in[172]), .N271(in[173]), .N274(in[174]), .N277(in[175]), 
.N280(in[176]), .N283(in[177]), .N286(in[178]), .N289(in[179]), 
.N293(in[180]), .N296(in[181]), .N299(in[182]), .N303(in[183]), 
.N307(in[184]), .N310(in[185]), .N313(in[186]), .N316(in[187]), 
.N319(in[188]), .N322(in[189]), .N325(in[190]), .N328(in[191]), 
.N331(in[192]), .N334(in[193]), .N337(in[194]), .N340(in[195]), 
.N343(in[196]), .N346(in[197]), .N349(in[198]), .N352(in[199]), 
.N355(in[200]), .N358(in[201]), .N361(in[202]), .N364(in[203]), 
.N367(in[204]), .N382(in[205]), .N241_I(in[206]), .N387(out[0]), .N388(out[1]), .N478(out[2]), .N482(out[3]), 
.N484(out[4]), .N486(out[5]), .N489(out[6]), .N492(out[7]), 
.N501(out[8]), .N505(out[9]), .N507(out[10]), .N509(out[11]), 
.N511(out[12]), .N513(out[13]), .N515(out[14]), .N517(out[15]), 
.N519(out[16]), .N535(out[17]), .N537(out[18]), .N539(out[19]), 
.N541(out[20]), .N543(out[21]), .N545(out[22]), .N547(out[23]), 
.N549(out[24]), .N551(out[25]), .N553(out[26]), .N556(out[27]), 
.N559(out[28]), .N561(out[29]), .N563(out[30]), .N565(out[31]), 
.N567(out[32]), .N569(out[33]), .N571(out[34]), .N573(out[35]), 
.N582(out[36]), .N643(out[37]), .N707(out[38]), .N813(out[39]), 
.N881(out[40]), .N882(out[41]), .N883(out[42]), .N884(out[43]), 
.N885(out[44]), .N889(out[45]), .N945(out[46]), .N1110(out[47]), 
.N1111(out[48]), .N1112(out[49]), .N1113(out[50]), .N1114(out[51]), 
.N1489(out[52]), .N1490(out[53]), .N1781(out[54]), .N10025(out[55]), 
.N10101(out[56]), .N10102(out[57]), .N10103(out[58]), .N10104(out[59]), 
.N10109(out[60]), .N10110(out[61]), .N10111(out[62]), .N10112(out[63]), 
.N10350(out[64]), .N10351(out[65]), .N10352(out[66]), .N10353(out[67]), 
.N10574(out[68]), .N10575(out[69]), .N10576(out[70]), .N10628(out[71]), 
.N10632(out[72]), .N10641(out[73]), .N10704(out[74]), .N10706(out[75]), 
.N10711(out[76]), .N10712(out[77]), .N10713(out[78]), .N10714(out[79]), 
.N10715(out[80]), .N10716(out[81]), .N10717(out[82]), .N10718(out[83]), 
.N10729(out[84]), .N10759(out[85]), .N10760(out[86]), .N10761(out[87]), 
.N10762(out[88]), .N10763(out[89]), .N10827(out[90]), .N10837(out[91]), 
.N10838(out[92]), .N10839(out[93]), .N10840(out[94]), .N10868(out[95]), 
.N10869(out[96]), .N10870(out[97]), .N10871(out[98]), .N10905(out[99]), 
.N10906(out[100]), .N10907(out[101]), .N10908(out[102]), .N11333(out[103]), 
.N11334(out[104]), .N11340(out[105]), .N11342(out[106]), .N241_O(out[107]));

initial begin
   $readmemb(INPUT_FILE, memory);

   f = $fopen(OUTPUT_FILE);

   for (i = 0; i < NUMBER_OF_TESTS; i = i+1) begin
      in = memory[i];
      #1;
      $fdisplay(f, "%b", out);
   end
   $fclose(f);
   $finish;
end

endmodule