module test_nor(N3, N2, N1);

input N1,N2;
output N3;


nor NOR2_1 (N3, N2, N1);
endmodule
